module part1 ( A, B, P );
  input [7:0] A;
  input [7:0] B;
  output [15:0] P;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391;

  INV_X1 U5 ( .A(A[4]), .ZN(n241) );
  NAND2_X1 U6 ( .A1(B[4]), .A2(A[3]), .ZN(n8) );
  NAND2_X1 U7 ( .A1(B[6]), .A2(A[0]), .ZN(n27) );
  NAND2_X1 U8 ( .A1(B[5]), .A2(A[1]), .ZN(n5) );
  XOR2_X1 U9 ( .A(n27), .B(n5), .Z(n71) );
  NAND3_X1 U10 ( .A1(A[2]), .A2(B[4]), .A3(n71), .ZN(n7) );
  INV_X1 U11 ( .A(A[0]), .ZN(n360) );
  INV_X1 U12 ( .A(B[5]), .ZN(n282) );
  NOR2_X1 U13 ( .A1(n360), .A2(n282), .ZN(n20) );
  INV_X1 U14 ( .A(n20), .ZN(n118) );
  NAND2_X1 U15 ( .A1(A[1]), .A2(B[4]), .ZN(n77) );
  NOR2_X1 U16 ( .A1(n118), .A2(n77), .ZN(n70) );
  OR2_X1 U17 ( .A1(A[2]), .A2(n71), .ZN(n6) );
  NAND2_X1 U18 ( .A1(n70), .A2(n6), .ZN(n9) );
  NAND3_X1 U19 ( .A1(n8), .A2(n7), .A3(n9), .ZN(n67) );
  NAND2_X1 U20 ( .A1(A[2]), .A2(n71), .ZN(n10) );
  NAND2_X1 U21 ( .A1(n10), .A2(n9), .ZN(n11) );
  NAND2_X1 U22 ( .A1(n11), .A2(A[3]), .ZN(n66) );
  NAND2_X1 U23 ( .A1(A[1]), .A2(B[6]), .ZN(n38) );
  NOR2_X1 U24 ( .A1(n20), .A2(n38), .ZN(n14) );
  NAND2_X1 U25 ( .A1(A[2]), .A2(B[5]), .ZN(n12) );
  INV_X1 U26 ( .A(B[7]), .ZN(n312) );
  NOR2_X1 U27 ( .A1(n312), .A2(n360), .ZN(n18) );
  XNOR2_X1 U28 ( .A(n12), .B(n18), .ZN(n13) );
  XNOR2_X1 U29 ( .A(n14), .B(n13), .ZN(n69) );
  NAND2_X1 U30 ( .A1(n66), .A2(n69), .ZN(n15) );
  NAND2_X1 U31 ( .A1(n67), .A2(n15), .ZN(n17) );
  NOR2_X1 U32 ( .A1(n241), .A2(n17), .ZN(n88) );
  NAND2_X1 U33 ( .A1(B[4]), .A2(A[4]), .ZN(n16) );
  AND2_X1 U34 ( .A1(n17), .A2(n16), .ZN(n89) );
  INV_X1 U35 ( .A(n38), .ZN(n21) );
  NOR2_X1 U36 ( .A1(n21), .A2(n18), .ZN(n19) );
  INV_X1 U37 ( .A(A[2]), .ZN(n123) );
  NOR3_X1 U38 ( .A1(n19), .A2(n282), .A3(n123), .ZN(n24) );
  NAND2_X1 U39 ( .A1(n21), .A2(n20), .ZN(n22) );
  NOR2_X1 U40 ( .A1(B[7]), .A2(n22), .ZN(n23) );
  NOR2_X1 U41 ( .A1(n24), .A2(n23), .ZN(n26) );
  INV_X1 U42 ( .A(A[3]), .ZN(n235) );
  OR2_X1 U43 ( .A1(n26), .A2(n235), .ZN(n35) );
  NAND2_X1 U44 ( .A1(A[3]), .A2(B[5]), .ZN(n25) );
  NAND2_X1 U45 ( .A1(n26), .A2(n25), .ZN(n37) );
  NAND2_X1 U46 ( .A1(n35), .A2(n37), .ZN(n30) );
  NAND3_X1 U47 ( .A1(n27), .A2(A[1]), .A3(B[7]), .ZN(n29) );
  NAND2_X1 U48 ( .A1(B[6]), .A2(A[2]), .ZN(n28) );
  XNOR2_X1 U49 ( .A(n29), .B(n28), .ZN(n34) );
  XNOR2_X1 U50 ( .A(n30), .B(n34), .ZN(n90) );
  NOR2_X1 U51 ( .A1(n89), .A2(n90), .ZN(n31) );
  NOR2_X1 U52 ( .A1(n88), .A2(n31), .ZN(n32) );
  INV_X1 U53 ( .A(A[5]), .ZN(n313) );
  NOR2_X1 U54 ( .A1(n32), .A2(n313), .ZN(n95) );
  NAND2_X1 U55 ( .A1(A[5]), .A2(B[4]), .ZN(n33) );
  AND2_X1 U56 ( .A1(n33), .A2(n32), .ZN(n96) );
  NAND2_X1 U57 ( .A1(n35), .A2(n34), .ZN(n36) );
  NAND2_X1 U58 ( .A1(n37), .A2(n36), .ZN(n61) );
  NOR2_X1 U59 ( .A1(A[0]), .A2(A[2]), .ZN(n39) );
  NOR3_X1 U60 ( .A1(n39), .A2(n312), .A3(n38), .ZN(n54) );
  NAND2_X1 U61 ( .A1(A[3]), .A2(n54), .ZN(n42) );
  INV_X1 U62 ( .A(B[6]), .ZN(n295) );
  NOR2_X1 U63 ( .A1(n295), .A2(n235), .ZN(n40) );
  NOR2_X1 U64 ( .A1(n54), .A2(n40), .ZN(n51) );
  INV_X1 U65 ( .A(n51), .ZN(n41) );
  NAND2_X1 U66 ( .A1(n42), .A2(n41), .ZN(n44) );
  NAND2_X1 U67 ( .A1(B[7]), .A2(A[2]), .ZN(n43) );
  XNOR2_X1 U68 ( .A(n44), .B(n43), .ZN(n46) );
  NAND2_X1 U69 ( .A1(A[4]), .A2(B[5]), .ZN(n45) );
  NAND2_X1 U70 ( .A1(n46), .A2(n45), .ZN(n63) );
  OR3_X1 U71 ( .A1(n241), .A2(n282), .A3(n46), .ZN(n60) );
  NAND2_X1 U72 ( .A1(n63), .A2(n60), .ZN(n47) );
  XNOR2_X1 U73 ( .A(n61), .B(n47), .ZN(n97) );
  NOR2_X1 U74 ( .A1(n96), .A2(n97), .ZN(n48) );
  NOR2_X1 U75 ( .A1(n95), .A2(n48), .ZN(n50) );
  INV_X1 U76 ( .A(A[6]), .ZN(n318) );
  OR2_X1 U77 ( .A1(n50), .A2(n318), .ZN(n150) );
  NAND2_X1 U78 ( .A1(A[6]), .A2(B[4]), .ZN(n49) );
  NAND2_X1 U79 ( .A1(n50), .A2(n49), .ZN(n152) );
  NAND2_X1 U80 ( .A1(n150), .A2(n152), .ZN(n65) );
  NOR3_X1 U81 ( .A1(n51), .A2(n123), .A3(n312), .ZN(n53) );
  NOR2_X1 U82 ( .A1(n235), .A2(n312), .ZN(n52) );
  NOR2_X1 U83 ( .A1(n53), .A2(n52), .ZN(n159) );
  NOR2_X1 U84 ( .A1(n54), .A2(n53), .ZN(n55) );
  NOR2_X1 U85 ( .A1(n235), .A2(n55), .ZN(n160) );
  OR2_X1 U86 ( .A1(n159), .A2(n160), .ZN(n57) );
  NAND2_X1 U87 ( .A1(A[4]), .A2(B[6]), .ZN(n56) );
  XNOR2_X1 U88 ( .A(n57), .B(n56), .ZN(n59) );
  OR3_X1 U89 ( .A1(n313), .A2(n59), .A3(n282), .ZN(n155) );
  NAND2_X1 U90 ( .A1(A[5]), .A2(B[5]), .ZN(n58) );
  NAND2_X1 U91 ( .A1(n59), .A2(n58), .ZN(n158) );
  NAND2_X1 U92 ( .A1(n155), .A2(n158), .ZN(n64) );
  NAND2_X1 U93 ( .A1(n61), .A2(n60), .ZN(n62) );
  NAND2_X1 U94 ( .A1(n63), .A2(n62), .ZN(n156) );
  XNOR2_X1 U95 ( .A(n64), .B(n156), .ZN(n149) );
  XNOR2_X1 U96 ( .A(n65), .B(n149), .ZN(n145) );
  NAND2_X1 U97 ( .A1(n67), .A2(n66), .ZN(n68) );
  XOR2_X1 U98 ( .A(n69), .B(n68), .Z(n109) );
  XNOR2_X1 U99 ( .A(n71), .B(n70), .ZN(n73) );
  NAND2_X1 U100 ( .A1(A[2]), .A2(B[4]), .ZN(n72) );
  XNOR2_X1 U101 ( .A(n73), .B(n72), .ZN(n81) );
  NAND2_X1 U102 ( .A1(A[3]), .A2(B[3]), .ZN(n74) );
  NAND2_X1 U103 ( .A1(n81), .A2(n74), .ZN(n114) );
  NAND2_X1 U104 ( .A1(A[2]), .A2(B[3]), .ZN(n117) );
  NOR2_X1 U105 ( .A1(n118), .A2(n117), .ZN(n80) );
  INV_X1 U106 ( .A(n117), .ZN(n76) );
  NAND2_X1 U107 ( .A1(A[0]), .A2(B[3]), .ZN(n232) );
  NOR2_X1 U108 ( .A1(B[5]), .A2(n232), .ZN(n75) );
  NOR2_X1 U109 ( .A1(n76), .A2(n75), .ZN(n78) );
  NOR2_X1 U110 ( .A1(n78), .A2(n77), .ZN(n79) );
  NOR2_X1 U111 ( .A1(n80), .A2(n79), .ZN(n116) );
  INV_X1 U112 ( .A(B[3]), .ZN(n184) );
  OR3_X1 U113 ( .A1(n235), .A2(n184), .A3(n81), .ZN(n113) );
  NAND2_X1 U114 ( .A1(n116), .A2(n113), .ZN(n82) );
  AND2_X1 U115 ( .A1(n114), .A2(n82), .ZN(n110) );
  NOR2_X1 U116 ( .A1(n109), .A2(n110), .ZN(n83) );
  NOR3_X1 U117 ( .A1(n83), .A2(n184), .A3(n241), .ZN(n85) );
  AND2_X1 U118 ( .A1(n109), .A2(n110), .ZN(n84) );
  NOR2_X1 U119 ( .A1(n85), .A2(n84), .ZN(n87) );
  NOR2_X1 U120 ( .A1(n87), .A2(n313), .ZN(n135) );
  NAND2_X1 U121 ( .A1(A[5]), .A2(B[3]), .ZN(n86) );
  AND2_X1 U122 ( .A1(n87), .A2(n86), .ZN(n136) );
  OR2_X1 U123 ( .A1(n89), .A2(n88), .ZN(n91) );
  XNOR2_X1 U124 ( .A(n91), .B(n90), .ZN(n137) );
  NOR2_X1 U125 ( .A1(n136), .A2(n137), .ZN(n92) );
  OR2_X1 U126 ( .A1(n135), .A2(n92), .ZN(n94) );
  NAND2_X1 U127 ( .A1(n94), .A2(A[6]), .ZN(n105) );
  NOR2_X1 U128 ( .A1(n318), .A2(n184), .ZN(n93) );
  NOR2_X1 U129 ( .A1(n94), .A2(n93), .ZN(n104) );
  OR2_X1 U130 ( .A1(n96), .A2(n95), .ZN(n98) );
  XNOR2_X1 U131 ( .A(n98), .B(n97), .ZN(n107) );
  OR2_X1 U132 ( .A1(n104), .A2(n107), .ZN(n99) );
  NAND2_X1 U133 ( .A1(n105), .A2(n99), .ZN(n102) );
  INV_X1 U134 ( .A(n102), .ZN(n101) );
  NAND2_X1 U135 ( .A1(A[7]), .A2(B[3]), .ZN(n100) );
  NAND2_X1 U136 ( .A1(n101), .A2(n100), .ZN(n148) );
  NAND2_X1 U137 ( .A1(n102), .A2(A[7]), .ZN(n146) );
  NAND2_X1 U138 ( .A1(n148), .A2(n146), .ZN(n103) );
  XOR2_X1 U139 ( .A(n145), .B(n103), .Z(n270) );
  INV_X1 U140 ( .A(n104), .ZN(n106) );
  NAND2_X1 U141 ( .A1(n106), .A2(n105), .ZN(n108) );
  XOR2_X1 U142 ( .A(n108), .B(n107), .Z(n260) );
  NAND2_X1 U143 ( .A1(A[4]), .A2(B[3]), .ZN(n112) );
  XNOR2_X1 U144 ( .A(n110), .B(n109), .ZN(n111) );
  XOR2_X1 U145 ( .A(n112), .B(n111), .Z(n133) );
  AND3_X1 U146 ( .A1(A[5]), .A2(n133), .A3(B[2]), .ZN(n203) );
  NAND2_X1 U147 ( .A1(n114), .A2(n113), .ZN(n115) );
  XOR2_X1 U148 ( .A(n116), .B(n115), .Z(n129) );
  AND3_X1 U149 ( .A1(n129), .A2(B[2]), .A3(A[4]), .ZN(n168) );
  XNOR2_X1 U150 ( .A(n118), .B(n117), .ZN(n120) );
  NAND3_X1 U151 ( .A1(B[4]), .A2(A[1]), .A3(n232), .ZN(n119) );
  XOR2_X1 U152 ( .A(n120), .B(n119), .Z(n127) );
  AND3_X1 U153 ( .A1(A[3]), .A2(B[2]), .A3(n127), .ZN(n192) );
  INV_X1 U154 ( .A(A[1]), .ZN(n383) );
  NOR2_X1 U155 ( .A1(n383), .A2(n184), .ZN(n173) );
  NAND3_X1 U156 ( .A1(A[0]), .A2(B[2]), .A3(n173), .ZN(n121) );
  NOR2_X1 U157 ( .A1(B[4]), .A2(n121), .ZN(n177) );
  INV_X1 U158 ( .A(B[4]), .ZN(n174) );
  NOR2_X1 U159 ( .A1(n360), .A2(n174), .ZN(n122) );
  NOR2_X1 U160 ( .A1(n173), .A2(n122), .ZN(n124) );
  INV_X1 U161 ( .A(B[2]), .ZN(n228) );
  NOR3_X1 U162 ( .A1(n124), .A2(n123), .A3(n228), .ZN(n125) );
  NOR2_X1 U163 ( .A1(n177), .A2(n125), .ZN(n194) );
  NOR2_X1 U164 ( .A1(n235), .A2(n228), .ZN(n126) );
  NOR2_X1 U165 ( .A1(n127), .A2(n126), .ZN(n193) );
  NOR2_X1 U166 ( .A1(n194), .A2(n193), .ZN(n128) );
  NOR2_X1 U167 ( .A1(n192), .A2(n128), .ZN(n170) );
  NOR2_X1 U168 ( .A1(n241), .A2(n228), .ZN(n130) );
  NOR2_X1 U169 ( .A1(n130), .A2(n129), .ZN(n169) );
  NOR2_X1 U170 ( .A1(n170), .A2(n169), .ZN(n131) );
  NOR2_X1 U171 ( .A1(n168), .A2(n131), .ZN(n205) );
  NOR2_X1 U172 ( .A1(n313), .A2(n228), .ZN(n132) );
  NOR2_X1 U173 ( .A1(n133), .A2(n132), .ZN(n202) );
  NOR2_X1 U174 ( .A1(n205), .A2(n202), .ZN(n134) );
  NOR2_X1 U175 ( .A1(n203), .A2(n134), .ZN(n211) );
  OR2_X1 U176 ( .A1(n136), .A2(n135), .ZN(n138) );
  XNOR2_X1 U177 ( .A(n138), .B(n137), .ZN(n210) );
  NAND2_X1 U178 ( .A1(n211), .A2(n210), .ZN(n141) );
  NAND2_X1 U179 ( .A1(A[6]), .A2(B[2]), .ZN(n212) );
  OR2_X1 U180 ( .A1(n210), .A2(n211), .ZN(n139) );
  NAND2_X1 U181 ( .A1(n212), .A2(n139), .ZN(n140) );
  AND2_X1 U182 ( .A1(n141), .A2(n140), .ZN(n259) );
  OR2_X1 U183 ( .A1(n260), .A2(n259), .ZN(n142) );
  NAND3_X1 U184 ( .A1(n142), .A2(A[7]), .A3(B[2]), .ZN(n144) );
  NAND2_X1 U185 ( .A1(n260), .A2(n259), .ZN(n143) );
  NAND2_X1 U186 ( .A1(n144), .A2(n143), .ZN(n269) );
  AND2_X1 U187 ( .A1(n270), .A2(n269), .ZN(n167) );
  NAND2_X1 U188 ( .A1(n146), .A2(n145), .ZN(n147) );
  NAND2_X1 U189 ( .A1(n148), .A2(n147), .ZN(n323) );
  NAND2_X1 U190 ( .A1(n150), .A2(n149), .ZN(n151) );
  NAND2_X1 U191 ( .A1(n152), .A2(n151), .ZN(n153) );
  INV_X1 U192 ( .A(A[7]), .ZN(n281) );
  OR2_X1 U193 ( .A1(n153), .A2(n281), .ZN(n305) );
  NAND2_X1 U194 ( .A1(A[7]), .A2(B[4]), .ZN(n154) );
  NAND2_X1 U195 ( .A1(n154), .A2(n153), .ZN(n307) );
  NAND2_X1 U196 ( .A1(n305), .A2(n307), .ZN(n165) );
  NAND2_X1 U197 ( .A1(n156), .A2(n155), .ZN(n157) );
  NAND2_X1 U198 ( .A1(n158), .A2(n157), .ZN(n286) );
  NAND2_X1 U199 ( .A1(B[6]), .A2(A[5]), .ZN(n162) );
  NOR2_X1 U200 ( .A1(n312), .A2(n241), .ZN(n294) );
  NOR3_X1 U201 ( .A1(n159), .A2(n295), .A3(n241), .ZN(n297) );
  NOR2_X1 U202 ( .A1(n297), .A2(n160), .ZN(n292) );
  XOR2_X1 U203 ( .A(n294), .B(n292), .Z(n161) );
  XNOR2_X1 U204 ( .A(n162), .B(n161), .ZN(n287) );
  XNOR2_X1 U205 ( .A(n286), .B(n287), .ZN(n164) );
  NAND2_X1 U206 ( .A1(A[6]), .A2(B[5]), .ZN(n163) );
  XNOR2_X1 U207 ( .A(n164), .B(n163), .ZN(n304) );
  XNOR2_X1 U208 ( .A(n165), .B(n304), .ZN(n322) );
  XOR2_X1 U209 ( .A(n323), .B(n322), .Z(n166) );
  NAND2_X1 U210 ( .A1(n167), .A2(n166), .ZN(n328) );
  OR2_X1 U211 ( .A1(n167), .A2(n166), .ZN(n327) );
  NAND2_X1 U212 ( .A1(n328), .A2(n327), .ZN(n274) );
  INV_X1 U213 ( .A(B[1]), .ZN(n384) );
  NOR2_X1 U214 ( .A1(n318), .A2(n384), .ZN(n200) );
  OR2_X1 U215 ( .A1(n169), .A2(n168), .ZN(n171) );
  XNOR2_X1 U216 ( .A(n171), .B(n170), .ZN(n198) );
  OR3_X1 U217 ( .A1(n313), .A2(n384), .A3(n198), .ZN(n215) );
  NOR2_X1 U218 ( .A1(n241), .A2(n384), .ZN(n190) );
  NAND2_X1 U219 ( .A1(A[2]), .A2(B[2]), .ZN(n181) );
  NAND3_X1 U220 ( .A1(n228), .A2(A[0]), .A3(B[4]), .ZN(n172) );
  NAND2_X1 U221 ( .A1(n172), .A2(n173), .ZN(n176) );
  OR3_X1 U222 ( .A1(n174), .A2(n360), .A3(n173), .ZN(n175) );
  NAND2_X1 U223 ( .A1(n176), .A2(n175), .ZN(n179) );
  INV_X1 U224 ( .A(n177), .ZN(n178) );
  NAND2_X1 U225 ( .A1(n179), .A2(n178), .ZN(n180) );
  XNOR2_X1 U226 ( .A(n181), .B(n180), .ZN(n187) );
  OR3_X1 U227 ( .A1(n235), .A2(n384), .A3(n187), .ZN(n237) );
  NAND2_X1 U228 ( .A1(A[1]), .A2(B[2]), .ZN(n182) );
  NAND2_X1 U229 ( .A1(n232), .A2(n182), .ZN(n183) );
  NAND3_X1 U230 ( .A1(n183), .A2(A[2]), .A3(B[1]), .ZN(n186) );
  NOR2_X1 U231 ( .A1(n360), .A2(n384), .ZN(n390) );
  NAND4_X1 U232 ( .A1(A[1]), .A2(B[2]), .A3(n390), .A4(n184), .ZN(n185) );
  NAND2_X1 U233 ( .A1(n186), .A2(n185), .ZN(n239) );
  NAND2_X1 U234 ( .A1(A[3]), .A2(B[1]), .ZN(n188) );
  NAND2_X1 U235 ( .A1(n188), .A2(n187), .ZN(n238) );
  NAND2_X1 U236 ( .A1(n239), .A2(n238), .ZN(n189) );
  NAND2_X1 U237 ( .A1(n237), .A2(n189), .ZN(n191) );
  NOR2_X1 U238 ( .A1(n190), .A2(n191), .ZN(n219) );
  AND2_X1 U239 ( .A1(A[4]), .A2(n191), .ZN(n220) );
  OR2_X1 U240 ( .A1(n193), .A2(n192), .ZN(n195) );
  XOR2_X1 U241 ( .A(n195), .B(n194), .Z(n221) );
  NOR2_X1 U242 ( .A1(n220), .A2(n221), .ZN(n196) );
  NOR2_X1 U243 ( .A1(n219), .A2(n196), .ZN(n218) );
  NAND2_X1 U244 ( .A1(A[5]), .A2(B[1]), .ZN(n197) );
  NAND2_X1 U245 ( .A1(n198), .A2(n197), .ZN(n216) );
  NAND2_X1 U246 ( .A1(n218), .A2(n216), .ZN(n199) );
  NAND2_X1 U247 ( .A1(n215), .A2(n199), .ZN(n201) );
  NOR2_X1 U248 ( .A1(n200), .A2(n201), .ZN(n251) );
  AND2_X1 U249 ( .A1(A[6]), .A2(n201), .ZN(n252) );
  OR2_X1 U250 ( .A1(n203), .A2(n202), .ZN(n204) );
  XOR2_X1 U251 ( .A(n205), .B(n204), .Z(n253) );
  NOR2_X1 U252 ( .A1(n252), .A2(n253), .ZN(n206) );
  NOR2_X1 U253 ( .A1(n251), .A2(n206), .ZN(n209) );
  INV_X1 U254 ( .A(n209), .ZN(n208) );
  NAND2_X1 U255 ( .A1(A[7]), .A2(B[1]), .ZN(n207) );
  NAND2_X1 U256 ( .A1(n208), .A2(n207), .ZN(n263) );
  NAND2_X1 U257 ( .A1(n209), .A2(A[7]), .ZN(n266) );
  NAND2_X1 U258 ( .A1(n263), .A2(n266), .ZN(n214) );
  XOR2_X1 U259 ( .A(n211), .B(n210), .Z(n213) );
  XNOR2_X1 U260 ( .A(n213), .B(n212), .ZN(n264) );
  XNOR2_X1 U261 ( .A(n214), .B(n264), .ZN(n374) );
  NAND2_X1 U262 ( .A1(n216), .A2(n215), .ZN(n217) );
  XOR2_X1 U263 ( .A(n218), .B(n217), .Z(n249) );
  INV_X1 U264 ( .A(B[0]), .ZN(n359) );
  OR3_X1 U265 ( .A1(n318), .A2(n249), .A3(n359), .ZN(n375) );
  OR2_X1 U266 ( .A1(n220), .A2(n219), .ZN(n222) );
  XOR2_X1 U267 ( .A(n222), .B(n221), .Z(n246) );
  OR3_X1 U268 ( .A1(n359), .A2(n313), .A3(n246), .ZN(n365) );
  NAND2_X1 U269 ( .A1(B[2]), .A2(A[0]), .ZN(n387) );
  NAND2_X1 U270 ( .A1(B[1]), .A2(A[1]), .ZN(n223) );
  NAND2_X1 U271 ( .A1(n387), .A2(n223), .ZN(n224) );
  NAND3_X1 U272 ( .A1(n224), .A2(A[2]), .A3(B[0]), .ZN(n227) );
  NAND2_X1 U273 ( .A1(A[1]), .A2(n390), .ZN(n225) );
  NOR2_X1 U274 ( .A1(n359), .A2(n225), .ZN(n385) );
  NAND2_X1 U275 ( .A1(n385), .A2(n387), .ZN(n226) );
  NAND2_X1 U276 ( .A1(n227), .A2(n226), .ZN(n371) );
  OR3_X1 U277 ( .A1(n390), .A2(n228), .A3(n383), .ZN(n230) );
  NAND2_X1 U278 ( .A1(A[2]), .A2(B[1]), .ZN(n229) );
  XNOR2_X1 U279 ( .A(n230), .B(n229), .ZN(n231) );
  XNOR2_X1 U280 ( .A(n232), .B(n231), .ZN(n234) );
  NAND2_X1 U281 ( .A1(A[3]), .A2(B[0]), .ZN(n233) );
  NAND2_X1 U282 ( .A1(n234), .A2(n233), .ZN(n369) );
  NAND2_X1 U283 ( .A1(n371), .A2(n369), .ZN(n236) );
  OR3_X1 U284 ( .A1(n235), .A2(n359), .A3(n234), .ZN(n370) );
  AND2_X1 U285 ( .A1(n236), .A2(n370), .ZN(n243) );
  NAND2_X1 U286 ( .A1(n238), .A2(n237), .ZN(n240) );
  XOR2_X1 U287 ( .A(n240), .B(n239), .Z(n242) );
  AND2_X1 U288 ( .A1(n243), .A2(n242), .ZN(n380) );
  NOR2_X1 U289 ( .A1(n241), .A2(n359), .ZN(n382) );
  NOR2_X1 U290 ( .A1(n243), .A2(n242), .ZN(n379) );
  NOR2_X1 U291 ( .A1(n382), .A2(n379), .ZN(n244) );
  NOR2_X1 U292 ( .A1(n380), .A2(n244), .ZN(n367) );
  NAND2_X1 U293 ( .A1(A[5]), .A2(B[0]), .ZN(n245) );
  NAND2_X1 U294 ( .A1(n246), .A2(n245), .ZN(n366) );
  NAND2_X1 U295 ( .A1(n367), .A2(n366), .ZN(n247) );
  NAND2_X1 U296 ( .A1(n365), .A2(n247), .ZN(n377) );
  NAND2_X1 U297 ( .A1(A[6]), .A2(B[0]), .ZN(n248) );
  NAND2_X1 U298 ( .A1(n249), .A2(n248), .ZN(n376) );
  NAND2_X1 U299 ( .A1(n377), .A2(n376), .ZN(n250) );
  NAND2_X1 U300 ( .A1(n375), .A2(n250), .ZN(n255) );
  NAND2_X1 U301 ( .A1(n255), .A2(A[7]), .ZN(n361) );
  OR2_X1 U302 ( .A1(n252), .A2(n251), .ZN(n254) );
  XNOR2_X1 U303 ( .A(n254), .B(n253), .ZN(n363) );
  INV_X1 U304 ( .A(n255), .ZN(n257) );
  NAND2_X1 U305 ( .A1(A[7]), .A2(B[0]), .ZN(n256) );
  NAND2_X1 U306 ( .A1(n257), .A2(n256), .ZN(n362) );
  NAND2_X1 U307 ( .A1(n363), .A2(n362), .ZN(n258) );
  NAND2_X1 U308 ( .A1(n361), .A2(n258), .ZN(n373) );
  NAND2_X1 U309 ( .A1(n374), .A2(n373), .ZN(n280) );
  XOR2_X1 U310 ( .A(n260), .B(n259), .Z(n262) );
  NAND2_X1 U311 ( .A1(A[7]), .A2(B[2]), .ZN(n261) );
  XNOR2_X1 U312 ( .A(n262), .B(n261), .ZN(n268) );
  NAND2_X1 U313 ( .A1(n264), .A2(n263), .ZN(n265) );
  NAND2_X1 U314 ( .A1(n266), .A2(n265), .ZN(n267) );
  XNOR2_X1 U315 ( .A(n268), .B(n267), .ZN(n279) );
  NOR2_X1 U316 ( .A1(n280), .A2(n279), .ZN(n277) );
  AND2_X1 U317 ( .A1(n268), .A2(n267), .ZN(n272) );
  XOR2_X1 U318 ( .A(n270), .B(n269), .Z(n271) );
  OR2_X1 U319 ( .A1(n272), .A2(n271), .ZN(n275) );
  NAND2_X1 U320 ( .A1(n277), .A2(n275), .ZN(n273) );
  NAND2_X1 U321 ( .A1(n272), .A2(n271), .ZN(n276) );
  NAND2_X1 U322 ( .A1(n273), .A2(n276), .ZN(n326) );
  XNOR2_X1 U323 ( .A(n274), .B(n326), .ZN(P[11]) );
  NAND2_X1 U324 ( .A1(n276), .A2(n275), .ZN(n278) );
  XNOR2_X1 U325 ( .A(n278), .B(n277), .ZN(P[10]) );
  XOR2_X1 U326 ( .A(n280), .B(n279), .Z(P[9]) );
  NOR2_X1 U327 ( .A1(n281), .A2(n282), .ZN(n289) );
  NOR3_X1 U328 ( .A1(n318), .A2(n282), .A3(n287), .ZN(n285) );
  AND2_X1 U329 ( .A1(n318), .A2(n287), .ZN(n283) );
  NOR2_X1 U330 ( .A1(n286), .A2(n283), .ZN(n284) );
  OR3_X1 U331 ( .A1(n289), .A2(n285), .A3(n284), .ZN(n308) );
  NAND2_X1 U332 ( .A1(n286), .A2(n318), .ZN(n291) );
  NAND2_X1 U333 ( .A1(n286), .A2(n287), .ZN(n290) );
  NAND2_X1 U334 ( .A1(n287), .A2(n318), .ZN(n288) );
  NAND4_X1 U335 ( .A1(n291), .A2(n290), .A3(n289), .A4(n288), .ZN(n311) );
  NAND2_X1 U336 ( .A1(n308), .A2(n311), .ZN(n303) );
  NAND2_X1 U337 ( .A1(B[7]), .A2(A[5]), .ZN(n302) );
  INV_X1 U338 ( .A(n292), .ZN(n293) );
  NOR2_X1 U339 ( .A1(n294), .A2(n293), .ZN(n296) );
  NOR3_X1 U340 ( .A1(n296), .A2(n295), .A3(n313), .ZN(n298) );
  NOR2_X1 U341 ( .A1(n298), .A2(n297), .ZN(n300) );
  NAND2_X1 U342 ( .A1(A[6]), .A2(B[6]), .ZN(n299) );
  AND2_X1 U343 ( .A1(n300), .A2(n299), .ZN(n314) );
  NOR2_X1 U344 ( .A1(n300), .A2(n318), .ZN(n315) );
  OR2_X1 U345 ( .A1(n314), .A2(n315), .ZN(n301) );
  XOR2_X1 U346 ( .A(n302), .B(n301), .Z(n309) );
  XOR2_X1 U347 ( .A(n303), .B(n309), .Z(n325) );
  NAND2_X1 U348 ( .A1(n305), .A2(n304), .ZN(n306) );
  NAND2_X1 U349 ( .A1(n307), .A2(n306), .ZN(n324) );
  NOR2_X1 U350 ( .A1(n325), .A2(n324), .ZN(n334) );
  NAND2_X1 U351 ( .A1(n309), .A2(n308), .ZN(n310) );
  NAND2_X1 U352 ( .A1(n311), .A2(n310), .ZN(n340) );
  NAND2_X1 U353 ( .A1(A[7]), .A2(B[6]), .ZN(n321) );
  NOR3_X1 U354 ( .A1(n314), .A2(n313), .A3(n312), .ZN(n316) );
  NOR2_X1 U355 ( .A1(n316), .A2(n315), .ZN(n319) );
  NAND2_X1 U356 ( .A1(A[6]), .A2(B[7]), .ZN(n317) );
  NAND2_X1 U357 ( .A1(n319), .A2(n317), .ZN(n336) );
  OR2_X1 U358 ( .A1(n319), .A2(n318), .ZN(n337) );
  NAND2_X1 U359 ( .A1(n336), .A2(n337), .ZN(n320) );
  XOR2_X1 U360 ( .A(n321), .B(n320), .Z(n341) );
  XOR2_X1 U361 ( .A(n340), .B(n341), .Z(n333) );
  NAND2_X1 U362 ( .A1(n334), .A2(n333), .ZN(n351) );
  NOR2_X1 U363 ( .A1(n323), .A2(n322), .ZN(n331) );
  XOR2_X1 U364 ( .A(n325), .B(n324), .Z(n330) );
  NAND2_X1 U365 ( .A1(n331), .A2(n330), .ZN(n355) );
  NAND2_X1 U366 ( .A1(n327), .A2(n326), .ZN(n329) );
  NAND2_X1 U367 ( .A1(n329), .A2(n328), .ZN(n357) );
  OR2_X1 U368 ( .A1(n331), .A2(n330), .ZN(n356) );
  NAND2_X1 U369 ( .A1(n357), .A2(n356), .ZN(n332) );
  NAND2_X1 U370 ( .A1(n355), .A2(n332), .ZN(n353) );
  OR2_X1 U371 ( .A1(n334), .A2(n333), .ZN(n352) );
  NAND2_X1 U372 ( .A1(n353), .A2(n352), .ZN(n335) );
  NAND2_X1 U373 ( .A1(n351), .A2(n335), .ZN(n349) );
  NAND3_X1 U374 ( .A1(n336), .A2(A[7]), .A3(B[6]), .ZN(n345) );
  NAND2_X1 U375 ( .A1(n345), .A2(n337), .ZN(n339) );
  NAND2_X1 U376 ( .A1(A[7]), .A2(B[7]), .ZN(n338) );
  XOR2_X1 U377 ( .A(n339), .B(n338), .Z(n342) );
  NAND2_X1 U378 ( .A1(n341), .A2(n340), .ZN(n343) );
  NAND2_X1 U379 ( .A1(n342), .A2(n343), .ZN(n348) );
  NAND2_X1 U380 ( .A1(n349), .A2(n348), .ZN(n346) );
  INV_X1 U381 ( .A(n343), .ZN(n344) );
  NAND4_X1 U382 ( .A1(B[7]), .A2(A[7]), .A3(n344), .A4(n345), .ZN(n347) );
  NAND3_X1 U383 ( .A1(n346), .A2(n345), .A3(n347), .ZN(P[15]) );
  NAND2_X1 U384 ( .A1(n348), .A2(n347), .ZN(n350) );
  XNOR2_X1 U385 ( .A(n350), .B(n349), .ZN(P[14]) );
  NAND2_X1 U386 ( .A1(n352), .A2(n351), .ZN(n354) );
  XNOR2_X1 U387 ( .A(n354), .B(n353), .ZN(P[13]) );
  NAND2_X1 U388 ( .A1(n356), .A2(n355), .ZN(n358) );
  XNOR2_X1 U389 ( .A(n358), .B(n357), .ZN(P[12]) );
  NOR2_X1 U390 ( .A1(n360), .A2(n359), .ZN(P[0]) );
  NAND2_X1 U391 ( .A1(n362), .A2(n361), .ZN(n364) );
  XNOR2_X1 U392 ( .A(n364), .B(n363), .ZN(P[7]) );
  NAND2_X1 U393 ( .A1(n366), .A2(n365), .ZN(n368) );
  XNOR2_X1 U394 ( .A(n368), .B(n367), .ZN(P[5]) );
  NAND2_X1 U395 ( .A1(n370), .A2(n369), .ZN(n372) );
  XNOR2_X1 U396 ( .A(n372), .B(n371), .ZN(P[3]) );
  XOR2_X1 U397 ( .A(n374), .B(n373), .Z(P[8]) );
  NAND2_X1 U398 ( .A1(n376), .A2(n375), .ZN(n378) );
  XNOR2_X1 U399 ( .A(n378), .B(n377), .ZN(P[6]) );
  NOR2_X1 U400 ( .A1(n380), .A2(n379), .ZN(n381) );
  XOR2_X1 U401 ( .A(n382), .B(n381), .Z(P[4]) );
  NOR3_X1 U402 ( .A1(n385), .A2(n384), .A3(n383), .ZN(n386) );
  XNOR2_X1 U403 ( .A(n387), .B(n386), .ZN(n389) );
  NAND2_X1 U404 ( .A1(A[2]), .A2(B[0]), .ZN(n388) );
  XNOR2_X1 U405 ( .A(n389), .B(n388), .ZN(P[2]) );
  NAND2_X1 U406 ( .A1(B[0]), .A2(A[1]), .ZN(n391) );
  XNOR2_X1 U407 ( .A(n391), .B(n390), .ZN(P[1]) );
endmodule

